/*
 Name: clk_gen.v
 Module: CLK_GENERATOR

 Output: CLK - output clock with period `SYS_CLK_FREQ

 Notes: Clock generator. The clock frequency is defined in the project definition file.
 

 Revision History:

 Version	Date		Who		email			note
------------------------------------------------------------------------------------------
  1.0     Sep 10, 2014	Kaushik Patra	kpatra@sjsu.edu		Initial creation
  2.0     Oct 29, 2014  David Thorpe    DE.Thorpe@gmail.com     Met output goals for DaVinci_TB
------------------------------------------------------------------------------------------*/
`include "prj_definition.v"
module CLK_GENERATOR(CLK);
    // output list;
    output CLK;

    // storage for clock value
    reg CLK;

    // Clock initialization
    initial begin
        CLK = 1'b1;
    end
    // For ever perform the following task.
    always begin
        #`SYS_CLK_HALF_PERIOD CLK <= ~CLK;
    end
endmodule
