`include "prj_definition.v"
/*
The gate based sequential multipler.
*/
module multiply(result, multiplicand, multiplier, write, shift, load);
	output [63:0] result;
	input [31:0] multiplicand, multiplier;
	input write, shift, load;
	wire [31:0] adderOut, andOut;
	wire dontCare;
	wire [63:0] shifterOut;

	reg [5:0] shiftNum;
	
	reg [63:0] result;
	reg [31:0] andProduct;

	and32 andGate(andOut, multiplicand, {32{result[0]}});
	rc_add_sub_32 adder(adderOut, dontCare, andOut, result[63:32], 1'b0);

	right_shifter64 b(shifterOut, result, shiftNum);

	initial shiftNum = {6'b000001};
	initial result = {{64'd0000},multiplier};
	
	always @(load) begin
		shiftNum = {6'b000001};
		result = {{64'd0000},multiplier};
	end
	always @(posedge write) begin
		result[63:32]=adderOut;
	end
	always @(posedge shift) begin
		result=shifterOut;
	end
endmodule
/*
The control unit for the sequential multiplier
*/
module mulControl(result, ready, multiplicand, multiplier, clk);
	output [63:0] result;
	output ready;

	input [31:0] multiplicand, multiplier;
	input clk;

	reg shift, write, load;
//unsignedWire[63:32], unsignedWire[31:0],
	mult mulPath(result[63:32], result[31:0], multiplicand,  multiplier, write, shift, load);

	reg [5:0] bit;
	wire ready = !bit;

	initial bit = 1'b0;
	initial load = 1'b1;
	always @( posedge clk )
		if(ready) begin
			bit = 6'b100000;
			load = 1'b0;
			write = 1'b0;
			shift = 1'b0;
		end else begin
			write = 1'b1;
			#1 shift = 1'b1;
			write = 1'b0;
			#1 shift = 1'b0;
 			bit = bit - 1'b1;
		end

endmodule
/*
Test Bench for sequential multiplier
Runs for the number of clock cycles required to complete multiplication
*/
module a_mul_TB;
	wire [63:0] result;
	wire ready;
	reg [31:0] multiplicand, multiplier;
	reg clk;

	mulControl mul(result, ready, multiplicand, multiplier, clk);

	initial begin
		multiplier = 32'b00010;
		multiplicand = 32'b0001;
		#1 clk = 1'b0; #1 clk = 1'b1; 
		#1 clk = 1'b0; #1 clk = 1'b1; 
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1; 
		#1 clk = 1'b0; #1 clk = 1'b1; 
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
		#1 clk = 1'b0; #1 clk = 1'b1;
	end
endmodule
module mult(resultHigh, resultLow, multiplicand, multiplier, write, shift, load);
	input [31:0] multiplicand, multiplier;
	output [31:0] resultHigh, resultLow;
	wire [31:0] bundle [3:0];
	wire [63:0] unsignedWire, twosOutm, muxOut;
	input write, shift, load;
	wire xorGate;

	xor o(xorGate, multiplicand[31], multiplier[31]);

	twosComplement t1(bundle[0], multiplicand);
	mux32_2x1 m1(bundle[1], multiplicand, bundle[0], multiplicand[31]);

	twosComplement t2(bundle[2], multiplier);
	mux32_2x1 m2(bundle[3], multiplier, bundle[2], multiplier[31]);

	//mult_32Bit_Unsigned mul(unsignedWire[63:32], unsignedWire[31:0], bundle[1], bundle[3]);
	multiply mulPath(unsignedWire, bundle[1], bundle[3], write, shift, load);

	twosComplement64 t3(twosOutm, unsignedWire);
	mux64_2x1 m3(muxOut, unsignedWire, twosOutm, xorGate);

	buf32 b1(resultLow, muxOut[31:0]);
	buf32 b2(resultHigh, muxOut[63:32]);
endmodule
